LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use IEEE.std_logic_unsigned.all;
 
ENTITY PC_tb IS
END PC_tb;
 
ARCHITECTURE behavior OF PC_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT PC
    PORT(
         CLK : IN  std_logic;
         rst : IN  std_logic;
         PCin : IN  std_logic_vector(5 downto 0);
         address : OUT  std_logic_vector(5 downto 0)
        );
    END COMPONENT;
    
   --Inputs
   signal CLK : std_logic := '0';
   signal rst : std_logic := '0';
   signal PCin : std_logic_vector(5 downto 0) := (others => '0');

 	--Outputs
   signal address : std_logic_vector(5 downto 0);

   -- Clock period definitions
   constant CLK_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: PC PORT MAP (
          CLK => CLK,
          rst => rst,
          PCin => PCin,
          address => address
        );

   -- Clock process definitions
   CLK_process :process
   begin
		CLK <= '0';
		wait for CLK_period/2;
		CLK <= '1';
		wait for CLK_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      wait for 100 ns;
		PCin <= address + '1';
      wait for 100 ns;
		PCin <= address + '1';
		rst <= '1';
      wait;
   end process;

END;
